PK   �"TT|$>�  �     cirkitFile.jsonݝYo#7ǿJ�}Uͻ�\���ͅ���GF�G���$� �}IY[�dw!��g���u���Xl5�/��n�n��n��;�m��ŕ�������Z?�m�\�nw��~��}���=�\�{�����~����]�5m����|Q��e[*�e�[S���՛��n����+l�4�v�.6ዲZv�uN��Z\/��g�x��g<�*�pW��-[Y��V�m]Q��4��TZ��׀g�5�`�Sw�z��{L]��	i�Kh��
�5�P�D\c�A��a2]W�8eWH���6mWlWzSץq�t���L
mP�6�l�UM���64��b�ڮ�˺i�~#M��?�l5���sk��M'��)��\�k�����^6�����!A���"���b�W�W��D	��^��K�{r����r 
�O��#������OR�>-t`���'��#�_�$���'��=I=��iؠ؁�	��ܒ��'@��D�E��ȶhq�O�q�o"���Md=4}������_��fe�uF��xo
ݖ}Q��cgZ/�N[����+�k�s�qj��vM��߹�	�t��Fӌ��:�q.T4=T�BU�BU�F���B��7
����O��i�?�A�4ȟ�3 �π���g@�ȟ�3 �ς�Y�?�珔��2&�Ο{�ML2�6�����Mz������%�܀?F\#�s�%��w�s>�?�A��fZN"<�I=�H���D< ��d>c#�EZ�&Lc�������6 �s�T�-q���C#�d7=�/p�&�X������$�� %��s�M�*A:�[Īĵ\\��x����`���oe��e���Z�D;��hj�b��Y�+�Ŋc�R�X�,V�	ވ.fF�ɲ��`ax����0��y<�e�c�D�����K�̙�Ͽv_#fx(�<K�8,y��X�P,y(V<+�c�)��X�P�f)�\1X��'j����Y�c1Xᙣ�@C��b�2f��Z�1��C���w>�#�tq��!X� <��˽8��P<��k�8��P<���8��P<���8̜(n*Ԍ8ә��Ȯ[Ν�uY��r�G*����)���P�x(V<+�X�xb��Ś'k�5SF�C��X�P�y(�<k�ņ�b�C���0�x(6<�ņ�b�C����Plg)�ց1Xs	$��j�-�J��O�ES��P��?�31����@��I�m�V)1X�]HԚ%�q�s�Q+zzd�V#��f�G��ѥ�L�,��(�=���L��Ld:2P+>>D��⍻c}���]w<�7`�nE�XQ,V4��bŲXq,V*+��:&xy�<�
~���`����aX�@,x(�<K��C��X�P,y(�<K�%Œ�b�C��X1�<+��,������<��7p+��D.������l�!o�Vf��x��:&xy�����fx �����fx�����Q������^��`������^��`������^��`������^��`�)��x>�o0��X�P�x(V<k�5Ś�b͔�P�y(�<k�5Ś�b�C����Plx(6L;�ņ�b�C����Ply(�<�Y�����ّ!o�Vx�2;I����l�!oLZ!o�Vf�\��[��#r�n�g�f�r�nev����V�������7p+���c�����{7����ŕ��ů�Cw������]ow������7�_�F��������|����:�V��/�k��R�w�rr��B�K�4qq@��^`���u��P�Ss��V]�Tu$��X�����2G$kG\#���eM��D�^�g��Q���Z�}��M�K_ ��P`me'��F��sM<M ��T_?�����}H��]���߄F~�d�::�5�5r���Jꎷ ��O-���|�b�@=J��$PO��5�RD�/6	�=��0$'�/���_p)�������c�:�?�1ȵ�U΃ �h4�X�蹔a��)���0�ao |fehzt�l�k�`��Y��yo|������ow��y��U����Eo��2�	����\&0���!�G��96ǀ��w�~�{P_�i�Zك��9�E�J���`A#n����EZ�L��}�@"�:�ޘ�B�K�b�^�F^�r*QN%ʩB9=�%��� J�BIT$��#�s@���O� �0����D  ��E�'� ��/� J�@�ʪ�wy!(��p*o��م�$N�M����ĩ̈~2��8��o�B�q�
{���U�W,�t�~%������B[z�-�a=
5�d)j�B���������Q05�l�$j�D���Q5J�FI4(�%Ѡ$�D�{PJ�AI4(�%Ѣ$Z�D��h'H$_ul��W��;���|�5�;��Ak2����_�:�D���~L��]XZ�G��i�:,�?���W`�C�Q$_���[��Xں%_��u�|_�6䋳s�!��`&2�%_��.�!7�N�uPȗk��x���̶�u��],d��F_\�YD�b���Ź��a���8��qN��zpdeE>�͝ʶD�QAD5N�D�j5dԐQCF5dԐQCE5ԩ9QCE/-(�_�K�?QCE5T��QCG5��QCG5t��QCG5L�0Q�Ds�t�0Q�D5L԰Q�F5l�q���O�(�[~>�J�����lB�4�(Kn��:����e��q���P07��W�u���������� ?�z2��meHF�Ճ�<��r<�Bd>�:{�$2��|%|�H��U�Ԏ�U@c�k����@c��O����q��i�9�r?w������m�5�-��hZ�������ԛ�&f.��Y�_���n�D���#u~�Ə���?��Gz�Ȝ��#{~dǏ���?�Ώ��#~�G���h��p��1����0����zs��v���u�_�l����9)���]��0훾!R�x&���[��?�æ�V뛮?F�2&���ﾪ�1W����o���p�v����]�_�)���x��~=�������r񾾹�?}~����n�,���������`wq��7w]xx�~��m77݇����o]��:���xW����9��M�|��=k�C�>CK�?+�����0o
Uʕ�Z:����T*ml�7m<�o���gt�y����p[�������p
?ֻ�A�t_.��m����e�������f{hn�󄾉���,�Y]����o
Y��~�t���ȳ��*'�Q�P-�K�*'W].'�ݜ��rJ\T��y���&����\��ܥ����Q�t9����P{a�܉�gra����h��he�he�����1[�1[i�\�1]�!^9�^�_�`i�1ai9᪕(/�=u��z|0�DdoS��ȍ�YM�7��>�_�����v�Sw�{�bU��Yt˭�'�ݶu��?�f��G����7 s��.Q��|����{�2a'uMQ�zS��w�������6�r�p�%�4�����x덡�b{u�����R7⌤f��7�z�m��+�ǒʮJ�$�UV�T#�ᤝZ�)�P��N\v�qWD�Iɤ��dڻ��=)����L{7侧$��S�i��=%����L{�OI���$�ޅ��=)����L{�.�Y����d�{J2��PG>))��S�b`��$��lfV���(rrv��S��I�"�L��II鲏�`���ލ۟����v����9Y��	�$\)�$[:L�ez�s�L�N�]���:!�v�L��j���|�$��S�I�ʓ��dz�NI����˒�i�)ɴw{�����Ӿ�iך��d�yJr���O�~�c!Tu�
��g�n��/�߱(�DK[9���L.��+[��c��o�'�v#��n��H�u8SU4U�k!�kO��	R��U������;~�c,�C��r&!�g��d8���I<4J.eH@*eT��Z+��S��{_���E�IUHe�N�emz14R��p�N���g0#�qL�2�,�^����e������4���|8��U�����|<c��~@�*i�=J�t6�1�ο��2t�	O�x�+m����z�Р��S��^�C���}d<�x8Y*��/�����}��B���J{�xW�z�T�D�=d����\)S�G>@
@i���;�G�G��19n)��O�2u.�J'�唠�D����D��!���ٛ)��aaZ�������M��]Ѻ���we�Z�u�z[���e=�(�h�ٿ��}|�s��؆gVjs0���~�8�1��ӄ�ο�i�-�}����|a˯�BV�}a�?��w�����e<;���*ē�7��T�)�Mf@�d؍E�Q��G�գݓT�H{�i�'$���N�sS��#�ղ"�5����PK   ܛ�SN��!I  I  /   images/bf4bccae-d76c-49e0-b144-227f603dc90a.png �@Y��PNG

   IHDR   p  	   L���   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  H�IDATx^�	�\U��_u���,$!Ye�]�QVqEG�9���Ց����u�st�`�7PT�î@�$l��H����������~շ��U��ם8��s��w����~w}���|�,N�0! �B��---A�X�A��#d2� ���l�=�}2ڸqc�y�{�S�;w��4������"l� ��-_�<Ȝz�Ž�޻���	F8�@&DL!(���A.�}�Ѡ���'��(ʹ#��E�"C%1������d50�X�vm"�at���Z|a툠"ԁ�a�W�`n ����Ą���QU+�#Ø�+�imo+�4�ie�[K�9����f�Z��j�`�W���ZبQ��ܴ.�	lk}�iy(*~�-sGE�.�I��l�[ۂ�lkP��KvkK6(�A6�nT6��#�O$L�y{3I�Z�	1�ݞac_ww�ߢ��ܵm۶�
��D���Z���Վ��?������=��
��f;�)BP��%���_\�y��Z�3f�Fu���GۦM�&�=~	�N&N�8Yᣣ,�{�, �6Ϙ�zh���իW��ꫯ.����c�y��#�xq��9���BO���[�n���=���~������c��Vy��ѣ'ϝ;wr�����<夓�x`ɓ�Np�"}���]�Y3�&�.&'���nԚ�ԪV�Qx�QG���3�|d�̙�/����r�nEj�U�Ώ?���;��~��}��w��F3�[(c3����G����M�=ۺ�3a ._��4���|P-��S� K06;#n$^&@�p��t7i��B�A�7�u��ocǎ�z����������~���Z1���	 �Z�ߴ%K������������:n�85��%>h:�ڣ!*@|0�	�z�FJl��h/1����?�9��`<��Įe��q�)/� ፂ�G%1���U�Vݲ뮻��E_|C[G���������+/����$�;�Lz\0,M�z�x���箮�~��4���&�|\�	��g�J�W� 2">ZA�4�� y�]��v�����޿�sν��̶(�!��]ӦM����^8o޼�k֬��0������B@�U�Ґ����E~�.�p��m�hǭ�!RF	A/nym��/��L�E�-Z�4a�sC�ҕ��(�BU�.MT�0{����>��{5ކM���m2Ǟ~��_�s�=�*�趶���@�a��7�=x���%P�����S��$�PQ7{���ߤ��Q�1z��n�Ur)nٲe[F���j1��'*p�{��.%� \��d�%@
��g�q�4�	���-�Q�������/|�F	EJ�]����;�w��sQH&Q>*@B3�`/]�D ޭ9����Q^�W��u�̓2kd(i,�aBtm�,Z%̌��"�ݵ`E0�AF#�7}�#Y6cƌ`¤�N�*�ר5�Z{��_s�w��&,�GީA��~�]w�w�%��s�����$��@H�"�2
�Fy��@
y�!�r��5�� �Bi��P��MP<C -�-��_^��ݍ�w]�*D����>�z-�׮[�x��0�Zvě\`� A�5��Y�i���$�i�/�(Ϯg�{��/��K�uZK�Ow�����֭[����b��hv-��aLx ���FZ� #0>n���U��b&�ڵkWt�A����1��o�r�)�,[�l�-@� ��M�����FȌ��a5��cK��h�xZ�p`:�$���Ν��}8$Z��w7(H���p�@���L��͐Wv�a/EQ�*��1k��ї^{����.�A �աs�hT�|�86t0ń��B�uu����2eʔ�.`���ٹYK��R"�R%��imLIތhT���.�g��$&0��K���CS�^-�^g,��A@��ֳ���@��\�&4�L�K���ݐ��.ʸ��FS4s7��2o�6*@�W��A ��3@�?Z�d{�=5�4���ѕ4�$�X���=h4$���9�ި�tO0�ঋ;�I�D��a��!�iiݺ�k,_��Su-�ZkB7��;d��m�B� �����"F�1p���t0ȴ��޼y���FG#0��Le�&�4�	��B"�CL�q��5jԬ�K���;�(��B>?��{�3qb��Lр	����k�<��X�$�w�yΝw޹��/4J�P,ZZ����~��ɓ'[��h4:Q6�o �#{�h��y��2F!03�}éS�N����zpH� ��ƽ�n�;�l�2���h��	�eSa�A-�������h��<k֬�����3L�B.�Q����?��[�Ν;���a��68��=0t�`�P�7��J�� �4��?������ԡ����/�|�]��=wƬ�%z�6��O� �>���0��^kh���d�h<�wk���foܸ�]+V�8T�#�%���Me�c����ʞL7l��[\e�1H�!��N�`���"l���X�h=�� �ɇu���g��?��O\���4̵jP�*���������7���sOW>��@O�CTf����ԍ�xV�O�M��ȴ���]{{{�Q�|̳H�,��͗{'��v��I2sdf)���2Z� 
��}�,�K��������O<��z��k��|�����K/���쳏���QXC^���N�>hrv��#����p���;*�9��-�������r!����/���dfѢE�'M��*��I��P�l��i"ԇ/�XT;��x�r��ӦMs���<�`��4o��4>��ѵ�����W�����nO�����zz[����ܙg�q��gϞEN�|���^,��K|�V��b�z���竴׊�`�l���;$�Gc���Hy �v�4ۓ�u��"2˜t�I�< s
�0�^�U�� B�i��\Z����ܖW��v�|0(Ųg�^%��㗿����~��>���'��ɶ��:�/��cW^}ձGu�$��ۺu�^�
h����^�a� }P��Ḝ�[�P���%'���ŷ���Γ��p�7?�/sq���7bg��")/u#��b�{��s�=�W�vح��yUh�h�[���<����iӦ��s�9�7n���'L�Vx@�9�����$�fӅB?��.���%�z��<�F ��Ȇ���8��8��I9�D�Bwv�`�hh*#D�T\�m[�t��u��-��׾v���X�_�Y�0��tqyȝU���Қm���ڵ�_���n���=��w�Y�KlX�?��=�z�Gx����s�"N�>h��1>��u=�Џ=�X�����kF _��L5A�1�@RH��'?��1��gzbʶ|�O _�u�]_8���"v�̙�uvv�g��!�{�i�>��'_2g˖-s�̙3z������ݿ³Sy;�V|:�h\ޢ��E�<�8r�8xM�-M�t�~��W�OS���'�R��#c��{�"��[a�e�P7Nd�SP��M9��m���h�����E?�ɏ�y睃��'t�2Im���	<�/��d[\���2{� /E�m<�l�q$y��@�y�.��Or��\�Qq�`�� �0�%"������(�Th��Z�k�#f�L,<�Ts�-Z�K�����pǀk�6�@i@�#�ܾQ6��s� G�Лzwp��U�n��u�C6����Gҍ�G��qf$<�p6F��E�Z0��g/����2"Z$bp�]
E���6XL&kl�<�HВ˅o�YS�m�����$�3<�mfKl���p�͇|��w_	�Τ4�)��9zϕ�Hxs�1�Ȇ�2���S� N7�i�'v���;�D$�%�1RZ���	O7�	����~?�Tຮ���=�	[�J+,�d"���Co#�D���0���i���E^� @��"ʸ>�	M�����e"�LG��GL$]+�pdD/)�aӦ ��v�<�I��[I�	Nݫ{%�����	O7 �&�vn7w�m��"}��m�Ე����2����t�	�8�@��������
*��LkeF��Gh&8�t���;*�X`��P	��Hx��@Z��dR�)�	O'�R6�lqK-�V�#>Tk`��$@�읩�j�	O7�G�xU'1�2	��ޑx����uy�xX�u`��!�, v�%t��,����LkeF�����u�v�z�Yn���0�����W���<��A'��IL���P�^	O?��dX�k��
ݲ�����:P�>%�H��u�����:��i�ׁ�YX��2#��W��bd����C��_9�f�����H[�F�k��C�:Ф\M����#�鄳���}d�� N>�����=��dX�kx�V�b�ԓ��l���;z8�ݧ��aH`���X���E��)�����f�aG7�l�"������50��m�����ϯ����cB��])<P�o����P��X/���p3�Z£��@�&����>߈c�|k�^x=��}p���%���Q��p	�?̍��x�?�y�l�,+�|C\��gp1��R����2�7B�e��D����Ƙ����4qy�u�e�?�>����∝	ƺRw��*0ar��*�KR~��j0��u �DM��֎u��]-����2}%����Z������~����S����0�w6δ��w`*¡�ʹf�Ѯ\�t���e�ۜ?yf�[z�\3��U��/�j��}ڻ�۽� �E����8:�Ϝ��׿z���s��{��^p�O/qژ)D���*.����}�q��w�Kӛ��ӧ�׭�=�G(e�*�y�;8��owq��������..���`��w.�����ѩJ*,������N��*��_�>8樣]���	&��ԙ�I'��2u:?5G�rº��;������~(�w�������O'�pB�ۂ!�e^��_���?��׾���ue��C>U�{�p��3�в�'nlhWG�h>�Â��p���E �L6��Kc��9�e��f�y�w�u�;�K8}�;�	~x��]� / 	��� |�%Ώ��!���o?�`�sχ��k�ҥ��I]EZ�8�������������7����J����wU)8%�R[���1��믿>�k�3���~o�$��,�e�u�Y�/o�9hS��k3*����7��m�.h'��7�tuu�}d���W�l��`����=�:������8" �ٺ-�m����?�x�5��:�&@�a�#�0���ҵ�)�0�Ry����;��9���Ki��k�`�D~Q-TZZ�*�M���\�j�*n����sP��o��˿���S	`ٲe��g�\y�.e(%�������&�2h}����$���,I�iӦ���.xe�jG-j�����^�[�,=�!�4&<W��+7e�B�!/���%}*$Pp5��2BK� ��)hbI�"�/?�i��XGc�Id��UW\��G���U:�T����l޼9���+]�SnQ<n� /��|����#\=¹��&*���a"'�O|��/��|�M�u��z�+�]y�߾�}�p��z�THY�J��O:�K=�t����L�y�+��s��V<�ܕ7o޼P������?���p
�������B���C�:���(#0&�9����zOh�1���.M��`ɒ%�to;�`w9�CJ]̒'��*��..�\l�կ~5����3���/���s����*;z��GE;�s��n��uo��C:�VJ��2��78׵�<wɺ��W�&N���h�(�=��#�o��z���B���;c<@ ��O�-빠8��]vY��,������o���o� ����v���EL��	�fKT֌K��F������� x��5�O�g���w_�u�n��a�c�y��`4��qcƸ2�}��/�	����_�]s��$̢�7��"-Z|�����w�uS�K+W���NY�L��� i�.yBs�0=��EcvVc��I�&�
)��=wn�m*.��g?��O
�z��~M|(���*u��i|�m��O_��̄�̱alI�^8O�A��T��:�֞|�	�Wei��~�d1��h��裏:7�)�2����2�T������'��\�d�B+c����o}����Z�׿�u�7ʳ⥕n�	H?g�G�1�.���~����-�<���7��Ёp�,�>��sխ������9>�����N�@�q�&�,a�n�#M5d�M<����Y�0�A�k�eL��Ø&��#K�ŋ��� c-��3Z�/7�  �5f ܹ��ҷ�4F1����?6H�0�^ �S�)�vv-@yb�nl~Ʌ_�����Ǝqy�t�1ʧkƏg�McǍsq��
Z;�<x�駃k��&X�b��-�ނ�<ݭ�A㥡��}h�� ��` �#.�.��[�"p�oݠ"�F�����T�a���a2�*��1@�V��.��}�jي�q$��O~�#���i�sI�`�?�x���?�я�Y'�#B��$���3N҂6-k������.?���|y�{�|���W���o�����v��q��~���ʻUJv�QG�<�'��|��*�#S	��E�	�g2wZ�BY$WN:���B7�b�'�t�H��λ�,�ō�Dˡǔ!�F ��&n�xLZ���M�=��#8T�+4�~�g���w�����h��g�q���a���6 0���̒�px�|xf���袋\�&�af����-9p[�FK-�]�	�fs���&�����j��I� �����u�b:���U⡇��)��q��kk���Z��3F(Rx��l7�(�	��)&n����$[]ĝ={���]�'���^r���E]�_�>��g6`��U�;G�?�l��)0WוFu�e�]�D�:�eU�~�9s��]�xQ>��ڃ������z�bm���UO>�H��)��M�8@�ς�R��}�s�����:�я~\|�������K.qS|N\j�W��7�J��=��C�������]��V1�4Ђ!3>Z.t���q��O�Jϖ�����d�q�:Q. S�ƍ�]z։��.Ӧ�PwG�r�׺�Z(t3�� ��ʗ�կ��f��^{��M [�lqt#x�l*�g�q��^�'�z([:!F��"-��d��@��F�t��GGsLp�;��ϻ5�zwp컎|�A��&Y�F�ݦn�w�}��T��ۺ\�_~\��>�M��'>eb�r��QnѮ�+F<���9�#d&$�*=kO��@�.��˂��������߃�O?ݵ�}��7����+/���A���O~\,��}ｎS�g%�M�t��wQ�4y���.�=�h��t�Y��m��U��[o���������?��@%�#��)3�Si���<�Ė@��V`�8�uuULV����Qb6��;\�#��-�$����o�t�Ť�{�ų���a:u��l8�d;(�Vw�f�Ld�R(h�ͯ~���_�6ٯ����]���^�<��}e������pՊ��W���_���������)���}�n՟�![}��n�g��Odǂ��B � ڹ#A�l�퓊�0F��
"�杕Ƒ��U���2��͛6�>��s����A|�Pl��V��k֬)�	C��Sn����Nsݚ��..��|~yp�7�|��_p���E8�䓃+���)�_&JFO��O<��cs�z�q@�~�?*2J)�Hq�ܦ'���;��j������
�� �7�fjQ���::{��.Q���S6��gh�o����	��'�Z�l�����c��|�>M��7f'�Қ����=[E�&-����m�&��9�Q�.�Z&6
�9zTеy�[�#|���S����>c�,�ۄ��W��1�V�c�/J!UV�h&݂��̙��q�&$��"�d�ۂ��QA�f�YjSZ&<�f�t���cluݻ¡��3~���F�Q��z`�uv���1d�w>ж��� �JUyUK-֒~����G�٠Z�~��ʼAe����?��gm��UY~ �i�!�7^��Z�Yxe����p?^s���WCe��&���۳o��ş8�)�G0��'��I�5Q�2	O7��ց����*6���^M>�s���|Ï8��u��P������/B�:���!	��]���
#�E�'&��J�0?�)[V�2��9	O7��m���s���=�ad����BQIGց���j��Gց;��3��«��]j��Z����eS���;^f�@�@�
$~�� |{����ʏ�R�M�4�X�3J����3I��|���/�l}˴V�`$<�p������k�"���!]PO�F0t@��ȷ�V,[$F|4�A`$���8��bׁDp���*0�\ib�#����7�a��3���_^n�vªA��q�S6��%�>��cWE�b�Ǵp��|x�W�?�>�
���j���}4�C�����"��M�i���,�����J�	ØnҸ�땗��@F�!ӌp���WӖ�0s����p��!�f�_3�aM|�_�Q�K��+��c�>�Z8�Ę<�m&�ٳ�|�LC�h��W�N���.���l	I�����b��8E��Q!��sx�W���yq��s��<a�B¢l��h �������]�CX����b�?w.����4.����Ew5���@a��0Sc�1aQ i�� �qGg�S�P�1�a7> ki	���a���)"�� o*ܧ��p�u���7�l.7G��4����`��
"�lԌU�;��� g8�ρN{�f2���Nl�plLN�r���dC*3_{l8G�������,����{c�:r=R81����Q�zձV���G�(O�΂=��>B�";��?�ض���"p���w�y������=:�Ł�"�1�����!@�Ќi�z���Q��\<�|��!V8l����v]w�����>�텓?����7*��st������s.�ܶ�>��_=���T�!��)oۖ.w����A��6�N�Ё�,z�e�R>�ih�qt'T�@�B mp]� !�[�&7�Z+ �w�y�ķg���L����r����P@�K�ٶNg�/���x{�Z���@B��,܄a=4��g�S(��8y4�g @�QD��$��]�j��縘�rd�`j��D�G�Nnܳz8E�.���9��h-0�p��ɒZ#)=K���4E�v�Š�����(G�1�Pȇ�$?hlo���૊���e�P3[	��Q}�>*8��?��a|�ćJ�,�C#��	37|e��%
�7���[�2��r�s�h���ΐ�Ɗ�Y���?���`�n�m�*4�gۃm��J��+ۮnNcWpP�U�ܕ��C&���+�j�����lu=�Y(��w�O;��S�k
Y弞+�I�mٜl&s���.�b���������J0mڴ�<��H�F�3�����؄k��U����yFa�
}X�?��9�Q�U�g����f�7Kt�$���)G�Gq��_������;>_�>
���[Z��O�
.Y@a�kgȡe!�4~�v��][�e	���?�Si8�v���\�X(~N���a�j���e {�on�m暫���w/�+��`T��i�،0�s�oy�[���O}K���
�R�Z�DU�����Ϲ���Rc5N�4�x�(�z�ʜ#s�7��Ε+W�;LSr'�UQ�$d|���<���@X��������*��_1=V�xCr�j��$ٓek��Mdo��Qv������e�.i���w�y�;S�5"m��#Hp��+I(�Ɋ��[dT� �k�}�m�bl��D�Mz�*�T!��2�x�-��^,{�]�cl���qV��T��=1e�
�9���!��������G�e��?��~^�2�˸i�Ei=���(�kf���d_#�Eiv�_.n�^��I�
�����?�~H�2�/�^/{���Uߧ��Z�_Q9��;�F�l���o���}nD�Wf�3z��jd6�,�9K��T�'4��l���[e��4����ܯ�v"���ge.U^N�	�_��L����2wȬQ�c+1��(h����\,�2��ߪa��ו7��]&��%U4 HYT������ "�м�d�;��H�h;����yJf�L�J�1����2w��.���A�[y\ ���c�L����A�>��ʄ��߫��� }�߃ `�&�SK�e�V��%D�Q\z��ո�K�<�	�?#��=� A�<3�i�{K��g�jϓ:��Hy�K���Oo�o������yT�� ��RО�]�av�ap*�����"3�fw�L��� ^���/l#���f�v������A�q��Wc#;���2;����%	��9�ltIp�I�/�|+Aq@����բܥ$�n� ?3vX8�3�(̖9Q嶱������OW%�N33��rR�����Kq4���-�z)ޮr��*PK��aợ:�N�
̰��R�n�Kc� �+d���	��U���Gl�Z��� ��!F��og��X/��������B�A-� ��7{4����1���� )�l����#���F:`��b�����Is('�d�
"Zʀ���f�gE\7_���]S����6!�X ��LM�|Th9И8� �[�Y��:������e2����v��E��Ҝ�P1��X@%}0�$��L�Ty���Rţ�S&v�QK��*��"��@��Ĕj�%���I#C��dx�X�h3%�(|��bi�%@C�ud�����	�v�9N�V=P&��3_h��Mc�TK�������bj��=9%f�����*�<$��1F11�ʊ���j��BWPly��'���I�{�U�� A�ߑ�{���K����%@(�dRĈ�Qאf�����m@�]�\��3�A��h��#�_\��0�d��U�u��
���
d�"���@��� �T�r`�*�e@}�W���j	�:
���l�И����E`�p�Lj4����k@��%�Z�Z$�� �d�๧����Js�T�&c|���;r3L��� �ց(J�+}�hT[���_%j
P&�-��,�������^+/t��I��e�Sp���H��� �f'�E��95QM3 &"h��)�Mseb5�inD#R6�����,�RP �Ίx�2l6����
P��|fE�$��7�R��<��Mh��2�՗�d�y���T��k2���h�yf0#�	L,�b��m�\�V-"� {f]#�=e�x�K�5������	lIq�bz���U���Z���.h`�i���A�'�����PK@H=�fB���qx�
�z5�W�{�J��'�%��i�@��b"�r���xg�o�B^&��8���[e`T���@���	�g�R��J�`O!(�����17���a�7�p��~VK��L���'�Q�
O�� ��˹�y�"���1�~�S�����1��q<�?��u�F����J"��*i��u�k�5C6�uY�{	*��|��*��>}�0l�q���gj	�.�n��P��� *� v�]ԝ1���R�Tr��ï"!�B�eH�o,�ʀe߆ք�->"B��V5ѧ�t-�ߛ�J�3g�˜&a�h�]�Ԣhf��ܱ�ki��F�i4}=��YE�h�Hhѓ�Dim�!���p�0VX7=zc{��z+�y�\s�m���o�6yr؅S �[���:��@9؉��?%�������N�J:�)��,T��w;�+_����¶�6���C:�8 Y��Y�M8k+�Y}�7�.���C=�-#��mm2T��K����ӿ���g���B!�i聏&,��D3��C#<�:����z�I�k����%�$��o��ڹ�,�X/�@�F���;��Ї
��r�A&���{�b0� ���׿~ٓO>���L�p�V�~���=,F�����a�9�c$@�6�!ٷ\{��G���`��E�#
��F.�����q���SO{\��q�ju�n���'�:u��t~��ֈ&a&N��?�=~�x�c�<�{�"��_��hyU4��3f�p��>}�������{�5k�s��&]p�q�tJ���7F��ҏ&�j��yڴ�ga�N�&�ND�h`�f-�~i��h�k6�ແ�(�V����6��H�y6?Z���ȬS�`�ʝ]����g3F����؆�}�S��Lb���a��0?��-���J����]��xc�=M���IEØ͆��<cx��0xV=��$�:��lgp�?@xfi���7��*�)@e\�"C
�P ���g�"�����d[[���H\Ҫ�h�`�Vj8ϑb�!�w���vz*i >O�v����3��cg�T�v�N� 3N�e��]�%��sw��k����|!O�݈mFKaF���yPi�1(��#�q�S`r&Hʻ��*J�0�Y� ]��4z�`\��v�x?����Y�Z=�u����4�� ��ȟ�� wRYn�C��=UҌ�3n3�y)]���/Q�a����[���˅A��F����+_R�m*+ؚ8��o#&\����p�"����5�*�R�h����=�Q>�j>�P�x�р/��Wf�M�zf/9��Q� ���`��&~�ABZ-�vU��|�*i�|6D4���J	��E��3��;<Ccߘ� �Õ���� ��^#�䫹Rj����;6���̀�+�M�t�1�2���r�)�Fc�HΰU8��<��Q?<`D�ML�d�>%�1��Yn}5�
&G����(��f�c����d������[d�^*�Z!��<�.,-R�ρ��6����hÖᖋ4'Y�!�� ]�>-F��gn�F�10v�+@e��m-�Z!	�. Ԏ�+�gB�P(Ν �� ���F��^����0/b+U���b��2����k=@��h���2�t�I(W��V���0��W�"�}�[�Z����Af*Q-�#���Ҽ��m��4���JB����i�i���$0|��g4z��֪� �����y9Ӗ���՝���5aQf١[�8�E�_����Ń�(��7��;@*�.PEw�gǠ�~Gc����|5�\p�.Y�M���[��Fk��BZY��4C���N��W�CUFk#��p�dd��~��2�>^�3�.4ZȻ�b��8z*O�QN.�I�R����2:���=y�`�[�D�8Z	A��+�°+�5�m�4��b�.U��>"��"A�-�����'�V?܇��ojbi�%@�F8G��}Qc ���A���U����`���CR��^}fߗ}>*������)m�U�� ���%�2��eh�Ռ����Ү?i��L _���8�m�|��(C�yߖ��r�ԣ�1��3�G#�����c��!��L+M��%��'Nhd���P�;!X ��e6=ЫF�O_=:�p�F_��T�1�?��J�)Gԅ2M�UF# z	�TA\���1ܽ�ȿ|�j�U�7ut������р�o`[iJS��^��-Ј��3 ��F@Z�
rK�J� z*�B���	��:���(�<��6����Z�颢w�;��0���a��#Z�a�Ms�%s�<�c���9��ҝ�,^��rŎQZQD���0��.f\�3C��@@X�������e�0�S�9�\�ʫ��JZ��"�p��JI�Sx�O�+i4�"��� ���8��F��ij8�Y�\���l2��Wk�զ*��� �P.e�:�~�uO�H�'�����F�RG��N�x�C����y�=^=&U���(LJ:���|�m�|��(C���}sQ�J�٧��q,�xbbyXK�4]�[�q%��
(�K����]�W����i\��l�o��E�� �C�-��� �u�`��&��7q��O`�S����¤F���Ȯ���4�1)j5��"z���=����	�	-zr A�D��16V��f�v�#��Ŧ�*@eF�Q۶���;+��ٰ;'c�'��#_βa�^$�ŗ���0M�G�[�.��V�jFZB�+7d��1a�#����"����Krw�)���t��ނ�	����C�a}K���O���/��K��Ζh%����-�s��	�d$>���,L!3�~���ǹ9F�♟@�{o1h�M��)O��w��Ȕ�F�-����p�k?K���&C�,fZZ֋?���l ���O�B��Ch�.D�?����*�*���իW��[���l
�+l���(�t�6o��}�ᦶ@�E��R�W��yES2 -&L��"�����[��̹GN��D��i�g˖��kk+��]�#���SxJn��o��� %��*y�����kgϞ���K/��H�`S�0l���-�|��/J{�TvUu�����?���g>�<G�)ߴ�}�c�J�f�W>�`���y*�D�z{z�����X@8��:;C��V�-�g�F�=�'r."v-K�
��Q�?9餓�������!�sC������6���V�Y_V6?S%R���1��v��5���0�e���Fx ��7O<�D��[nyRy|[a��a��
��|B�P8��#�|�;�:��^��a��z/�dn���=�\rɝ�g�:K�U=^bGeJ��=,�\{���s�=E����]s�T�f#<������x��	55��}мAϟ�������H�FZJ&�������q�,���ȴ8�B4}���/D(�� �!4 �&�\�bE�����7���b`��*~��w��u�M7��c`̡@���;����>ƏI�Xq��c��n������W�-Z<��3�.�&��Q�C��o|�k̘1+����6_	bN3�{f�:�{R�-K�.u�o�F�6I�k^}uÙ���74[� jM� PAyi�/�|Q��N�R�	�g���on���A��!��_��_'g�g�0^Cta�$@ρP.\���I�\�A�P�oN8�Ǹ�����a������Ţ��߭������*$G�0����
�'��RX��@�R���|�@�	a6�R�����<���kD����n�	]�g5��رc��-~����zH*@���p�[��d����2U�n-Dc��m�
/��!�:� ��=��+�\���2�8$ ���:���.��9�޿����v��i^+R�D�;in�O8>㫞�
���u�T��]��Y)���L�_yUET�Geb�n�����_��Ds4]���>��P��+��� ���LȻ���2�N�k�_��׺|&E�+8��j�`�UU,�[�P~|}�� w�I[ �lx5TV�
F�@��O@�|ǃv�
̖a�3�M���;iBū6�?�1X�%�[.� �W�YSIV�4�� ���v`�1 �ҹ�@��,r9\�I��l�>}� �)'~G�H�ʓ�S��_����L`��1�9e���)�Hh��r�.��{F&�_ $���Y�B����^KF�-*8Q�i���	v���1���۹���EJ�u���{L�a:S⣻�/�_K��ܦ��fo�a�:\�IZ~�V:�Qn�O��L
�W��K���{��3PQ8��aa�@���aS�P� &X���>D(��{��l	�Y|❢��{JRq
�I�Qv?����5��իG��z��ш e���p�L�vW ��ߥ��G�'<��C��P%��En��� ©��C��_�YK�X+�VZf,�^
�yB��0�\�Gj1Ɛ$Nڨ�dp�v�t����l��a��.�PK@���	ab��,��h4��������]^ч���*� �����M���c��y�]B>�@{�Z ���/��Ru���6e��U�S���)���I��>�XO2T��a�P��>Z_��|���$�X�C`"���؟�Db����ڢ�Q4\���;`�G��:�-��D���@�
�D��@Z`l\
���
m2��Ӭ����Pf��
֠���o�֨p93��\$ ��<L��i��4k�p��}����6�q�����2#��\�?� 4�~��`�J<�M�_o�B�~uJ�W��V����	��>��))V+��X&Ԣ���ݍr=w}��b$��K���6�cg�*�Y�ax� 9�_&@��1�����@uT�*�lc�.x�G↕(�
*�v���dzig|�Q����k�b⦯,�}�6��"�L@�#��t9^غu+�����ʫL��X���k]$ f���)V(���M� H�C��2E����o��	���s�����b��� eq��y4@ ���H`%����\v�1�I���$b�I��; �}ū~|7!�a���e���(R$,����� U0�@vb� yV�܈^���a� �MBB�c	� eQ�D�I*@2���]�� Mc �l6��;ɩ��ĭ� ���������������=%��>��g��^�D�I$@�Uύ�Á�<�P0�_�G}$Ұb�L=��(�P�i�{TvI8��L�S����V�����\.7���P�>F�ǲ�S�ԅ_b)���N�4zoKC� �GU@�O���pKO*�����PP�P�IڢAS�P�z�I���@��P����G�>�Q���%b����.`��4���M�DcdB�i@@���	� :�h����Z�-��]��}���0�� ���n�O�F�}@�1���7�oyd� }fx��c?A�a�7�.1ҧ/����!� �5���PN�
����z���[�FLq�=2���d��}�l'@�6��GW�%jI�U����j.-P� �T���W��Q�d��I��a���le�u�W�6�
�� p�h�� 
V��B�OR�.2}�ό��Q�����0V|t�[BO��� �I8���3�R��(T�`�H����U�a`8?��&��e�3��-���N&���,HH��	�a]h����cq����w%�ٻ�Z���g�E6��'eW����
P����\rDa���%��=���D��%bLJ� :�]�<���d��ԝw�f6��לL�
�jFkA��9�ba�����0�Nl~�2cRA��+��Iշ���s顕U
+f3�[�����DH$@�1�->+�%r97�9E����,�,yW=&>8�l�1�Z���xW�S�����J��E��(�
3�O��o�x/%@TY�=� ~�t�6�#�ۮ��"��d��9� Q��ʼ���#B],T��5 ˘�}�+u�l"!�>��郏� +Y"�6��M��PP��_�s��>,�������Do�T��b�M_���L��3!P���=ޣ����Y&m�|Ǹ3B2f��H^���|$�뤲:U���i��8A.�C��p��ͧ/�#=I�	P���~������}.7L��~����8��� 5ޕm�AAbG"�B�8K3�R�
�a�R?\`�B�����sd�E�L��̄�n�3�Et�g5�!� �7g��\�ʌ����{d�Zs�b�A�1ݢg�cЩĴ{�̰P<i���G����n����p�q]`$�
��%�0P0
sX|&���4 ��o���!Sh4Z����s��7,����֭[gJXN8(�E�sq"��EYW��c`Wwo��\��R(��m۶1=�E�P���N�0���0��l^�%�������WJ�9�
�s$��5/	PL(nذ!�oB<��S��O?�̒%K��?X�v-��w���$C1%#F���g��|ٲe���>������yY����s�;�������_��m�>�h�j�*~0A���zH��*��^|���o����m�hx&��Zb>_(�H���c�7-Z�S��I���!�hlW�������S�W��'k\��(Z>v��ࠃ��o�����3$DI��מ�ͷ�r˼ѣ;7�7�j��������p@硇z������_�' vWAm��� �˵�1Y�s���[��~����ĸ�����M�� ��zf^Q���������A�얆w��(��n_�^'�E߯�dC
��PYg������,��F�+'zr�J�������P}^����� ��|`��ӥ#�    IEND�B`�PK   �"Tx�H
c  �     jsons/user_defined.json��[k1����YC����}j)��R�d��m`M��TD��h�[���9�3��C~�K4A�I�Z�FiY�!���)��@0�^\��ԡ����q���{�`c��M�y+Kن�{c�)��5vF�]��.�!R5ث&���rT�B��R�QE�l�$�)HZ��p�Ą'��� �3ͤV�����^�+��-�z��1h�C:�g���NMC#�ZR�sii6�D&cJؑp�P��=@=��U��UF�q*]�^��4%�0Iq�Q��B�-ތ�iΎW2ʕ�G���xz�O�'�4~���.��܏����'�"a��d��M��V�E=/o���]QoM/�W���!���/ܯ��PK
   �"TT|$>�  �                   cirkitFile.jsonPK
   ܛ�SN��!I  I  /             �  images/bf4bccae-d76c-49e0-b144-227f603dc90a.pngPK
   �"Tx�H
c  �               $[  jsons/user_defined.jsonPK      �   �\    